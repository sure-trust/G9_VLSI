`timescale 1ns / 1ps
module decode4_16(y,a);
output reg [15:0]y; input [3:0]a;
always@(*) begin 
y[0]=(~a[3]&~a[2]&~a[1]&~a[0]);
y[1]=(~a[3]&~a[2]&~a[1]&a[0]);
y[2]=(~a[3]&~a[2]&a[1]&~a[0]);
y[3]=(~a[3]&~a[2]&a[1]&a[0]);
y[4]=(~a[3]&a[2]&~a[1]&~a[0]);
y[5]=(~a[3]&a[2]&~a[1]&a[0]);
y[6]=(~a[3]&a[2]&a[1]&~a[0]);
y[7]=(~a[3]&a[2]&a[1]&a[0]);
y[8]=(a[3]&~a[2]&~a[1]&~a[0]);
y[9]=(a[3]&~a[2]&~a[1]&a[0]);
y[10]=(a[3]&~a[2]&a[1]&~a[0]);
y[11]=(a[3]&~a[2]&a[1]&a[0]);
y[12]=(a[3]&a[2]&~a[1]&~a[0]);
y[13]=(a[3]&a[2]&~a[1]&a[0]);
y[14]=(a[3]&a[2]&a[1]&~a[0]);
y[15]=(a[3]&a[2]&a[1]&a[0]);
end
endmodule
