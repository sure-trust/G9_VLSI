`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:48:47 08/27/2023
// Design Name:   single_port_ram
// Module Name:   /home/student/Desktop/Sure Trust/RAM/single_port_ram_tb.v
// Project Name:  RAM
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: single_port_ram
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module single_port_ram_tb();

reg [7:0] data;
reg [5:0] address;
reg en,write_enable, clk;
wire [7:0] q;

single_port_ram dut(data, address, en,write_enable, clk, q);

initial begin
    clk=1'b1;
    forever #5 clk=~clk;
end

initial begin
    data= 8'h18;
    address= 6'd16;      
    en = 1'b1;write_enable= 1'b1;
    #100;
    
    data= 8'h29;
    address= 6'd12;      
    #100;
    
    data= 8'hAA;
    address= 6'd7;      
    #100;
	
	
    data= 8'hz; //read operation
    address= 6'd16;      
    write_enable= 1'b0;       
    #100;
    
    address= 6'd12;     
    #100;
    
    address= 6'd7;
    #100;
end

initial begin
$monitor("en: %b  write enable: %b  address: %d  data: %h  output: %h", en, write_enable, address, data, q);
#10000 $finish;
end
endmodule